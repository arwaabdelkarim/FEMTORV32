`timescale 1ns / 1ps
/******************************************************************* 
* 
* Module: Inst_Mem.v 
* Project: Arch_proj1 
* Author: Arwa Abdelkarim arwaabdelkarim@aucegypt.edu
          Farida Bey      farida.bey@aucegypt.edu
          
* Description: 
* 
* Change history: 
**********************************************************************/

module Inst_Mem(
    input [7:0] Addr,
    output [31:0] Data_out
    );
    
endmodule
